module decoder(inst_encoding, we);

input inst_encoding[31:0];
output we;





endmodule
